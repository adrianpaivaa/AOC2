library verilog;
use verilog.vl_types.all;
entity FULL_ADDER_1bit_vlg_sample_tst is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        CIN             : in     vl_logic;
        EN              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end FULL_ADDER_1bit_vlg_sample_tst;
