library verilog;
use verilog.vl_types.all;
entity REGISTER_BANK_vlg_vec_tst is
end REGISTER_BANK_vlg_vec_tst;
