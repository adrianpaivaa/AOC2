library verilog;
use verilog.vl_types.all;
entity DECODER_2X4_vlg_vec_tst is
end DECODER_2X4_vlg_vec_tst;
